.title KiCad schematic
.include "C:/AE/TLP290/tlp290_SE.mod"
XU1 /IN /K 0 /OUT TLP290_SE
R1 /OUT VDD {RC}
V2 VDD 0 DC {VSOURCE}
V1 /IN 0 sine({voff} {vampl} {freq})
R2 0 /K {RK}
.end
